//P176_七位显示译码器_74HC4511
module disp_decoder(
	input LE,BL,LT,	//LE,BL,LT为使能信号, LT,BL为低有效测试信号
	input [3:0] D,		//D为待显示的四位二进制数字
	output reg [6:0] L);   //L为7段显示器各段的工作情况

	wire [2:0] E;   
	assign E={LE,BL,LT}; //中间变量用于判断控制端优先级
	
	always@(*)
	begin
		 if(LE==0 && BL==1 && LT==1) 	//锁存器不工作
			begin		//译码器随输入变化
			  case(D)
				 //0-9显示。
				4'b0000:L=7'b111_1110;
				4'b0001:L=7'b011_0000;
				4'b0010:L=7'b110_1101;
				4'b0011:L=7'b111_1001;
				4'b0100:L=7'b011_0011;
				4'b0101:L=7'b101_1011;
				4'b0110:L=7'b001_1111;
				4'b0111:L=7'b111_0000;
				4'b1000:L=7'b111_1111;
				4'b1001:L=7'b111_1011;  
				//以下为无效状态
				4'b1010:L=7'b000_0000;
				4'b1011:L=7'b000_0000; 
				4'b1100:L=7'b000_0000;
				4'b1101:L=7'b000_0000;
				4'b1110:L=7'b000_0000;
				4'b1111:L=7'b000_0000; 		
				endcase
			end
		 else 
			begin
				casex(E)
				3'bxx0:L=7'b111_1111;  	//灯测试
				3'bx01:L=7'b000_0000; 	//灭灯
				3'b111:L<=L;				//锁存
				endcase
			end
	end
endmodule
